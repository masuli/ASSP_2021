module pc_init (zeros);

	parameter width = 0;

	output [width:0] zeros;
			
	assign zeros = 0;

endmodule 