package toplevel_imem_mau is
   -- created by generatebits
   constant IMEMMAUWIDTH : positive := 172;
end toplevel_imem_mau;
